// $Id: $
// File name:   Y_conv.sv
// Created:     12/2/2017
// Author:      Michael Karrs
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: Y Convolutionj Block.
