// $Id: $
// File name:   tb_image_buffer.sv
// Created:     12/4/2017
// Author:      Michael Karrs
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: Test Bench for Image Buffer.
